package common is
    constant INSTRUCTION_WIDTH: natural := 32;
end common;